<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-5.42907,11.7665,101.629,-42.025</PageViewport>
<gate>
<ID>2</ID>
<type>AA_FULLADDER_1BIT</type>
<position>32,-9.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_B_0</ID>26 </input>
<output>
<ID>OUT_0</ID>31 </output>
<input>
<ID>carry_in</ID>12 </input>
<output>
<ID>carry_out</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_FULLADDER_1BIT</type>
<position>43.5,-8.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_B_0</ID>24 </input>
<output>
<ID>OUT_0</ID>33 </output>
<input>
<ID>carry_in</ID>11 </input>
<output>
<ID>carry_out</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_FULLADDER_1BIT</type>
<position>56.5,-9.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_B_0</ID>5 </input>
<output>
<ID>OUT_0</ID>35 </output>
<input>
<ID>carry_in</ID>10 </input>
<output>
<ID>carry_out</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_FULLADDER_1BIT</type>
<position>71,-8.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_B_0</ID>3 </input>
<output>
<ID>OUT_0</ID>37 </output>
<input>
<ID>carry_in</ID>1 </input>
<output>
<ID>carry_out</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>10</ID>
<type>FF_GND</type>
<position>83.5,-10.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_MUX_2x1</type>
<position>21.5,-9.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>45 </output>
<input>
<ID>SEL_0</ID>100 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_FULLADDER_1BIT</type>
<position>34.5,-23.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_B_0</ID>26 </input>
<output>
<ID>OUT_0</ID>32 </output>
<input>
<ID>carry_in</ID>29 </input>
<output>
<ID>carry_out</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_FULLADDER_1BIT</type>
<position>47,-23.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_B_0</ID>24 </input>
<output>
<ID>OUT_0</ID>34 </output>
<input>
<ID>carry_in</ID>28 </input>
<output>
<ID>carry_out</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_FULLADDER_1BIT</type>
<position>59,-23.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_B_0</ID>5 </input>
<output>
<ID>OUT_0</ID>36 </output>
<input>
<ID>carry_in</ID>27 </input>
<output>
<ID>carry_out</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_FULLADDER_1BIT</type>
<position>72.5,-23.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_B_0</ID>3 </input>
<output>
<ID>OUT_0</ID>38 </output>
<input>
<ID>carry_in</ID>101 </input>
<output>
<ID>carry_out</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>239</ID>
<type>AA_TOGGLE</type>
<position>28,2.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_TOGGLE</type>
<position>35.5,2.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>241</ID>
<type>AA_TOGGLE</type>
<position>40.5,2.5</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>242</ID>
<type>AA_TOGGLE</type>
<position>46.5,2.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_MUX_2x1</type>
<position>34.5,-28.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>41 </output>
<input>
<ID>SEL_0</ID>100 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>243</ID>
<type>AA_TOGGLE</type>
<position>53,3</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_MUX_2x1</type>
<position>49,-29.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>42 </output>
<input>
<ID>SEL_0</ID>100 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>244</ID>
<type>AA_TOGGLE</type>
<position>60,2.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_MUX_2x1</type>
<position>63,-30</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>43 </output>
<input>
<ID>SEL_0</ID>100 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>245</ID>
<type>AA_TOGGLE</type>
<position>66,2.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_MUX_2x1</type>
<position>75.5,-29.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>44 </output>
<input>
<ID>SEL_0</ID>100 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>246</ID>
<type>AA_TOGGLE</type>
<position>73.5,3.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>36,-37.5</position>
<input>
<ID>N_in3</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>GA_LED</type>
<position>50,-38</position>
<input>
<ID>N_in3</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>254</ID>
<type>AA_TOGGLE</type>
<position>89.5,-29.5</position>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>63</ID>
<type>GA_LED</type>
<position>64.5,-38</position>
<input>
<ID>N_in3</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>256</ID>
<type>EE_VDD</type>
<position>79.5,-21.5</position>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>65</ID>
<type>GA_LED</type>
<position>76,-38</position>
<input>
<ID>N_in3</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>GA_LED</type>
<position>12.5,-10</position>
<input>
<ID>N_in1</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>48.5,11</position>
<gparam>LABEL_TEXT Carry Select Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>66,4.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>73,5.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>53,5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>40.5,5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>27.5,5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>60,4.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>46.5,4.5</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>35,5</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AA_LABEL</type>
<position>32.5,-19</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>35.5,-19</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>44.5,-19</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>49,-19.5</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>57.5,-19</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>60.5,-18.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>70,-19</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>73.5,-19</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_LABEL</type>
<position>81.5,-7</position>
<gparam>LABEL_TEXT Asumming Cin=0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_LABEL</type>
<position>83,-19</position>
<gparam>LABEL_TEXT Asumming Cin=1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>76,-41</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>64,-40.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>50,-40.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>35.5,-41</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>AA_LABEL</type>
<position>6,-10</position>
<gparam>LABEL_TEXT Cout</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>AA_LABEL</type>
<position>89,-26.5</position>
<gparam>LABEL_TEXT Select</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>32.5,-4.5</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>43,-4.5</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>56,-5.5</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>70,-4</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>72,-17</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>58.5,-17</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>AA_LABEL</type>
<position>47,-17</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>34,-16.5</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AA_LABEL</type>
<position>34.5,-31</position>
<gparam>LABEL_TEXT 2:1 MUX</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>AA_LABEL</type>
<position>49,-32</position>
<gparam>LABEL_TEXT 2:1 MUX</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>64,-32.5</position>
<gparam>LABEL_TEXT 2:1 MUX</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>76,-32.5</position>
<gparam>LABEL_TEXT 2:1 MUX</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>22,-13</position>
<gparam>LABEL_TEXT 2:1 MUX</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-8.5,83.5,-8.5</points>
<connection>
<GID>8</GID>
<name>carry_in</name></connection>
<intersection>83.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83.5,-9.5,83.5,-8.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-1,73.5,1.5</points>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>-1 3</intersection>
<intersection>0 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>72,-1,73.5,-1</points>
<intersection>72 4</intersection>
<intersection>73.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>72,-5.5,72,-1</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-1 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>73.5,0,76.5,0</points>
<intersection>73.5 0</intersection>
<intersection>76.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>76.5,-20.5,76.5,0</points>
<intersection>-20.5 8</intersection>
<intersection>0 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>73.5,-20.5,76.5,-20.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>76.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-5.5,70,-1.5</points>
<connection>
<GID>8</GID>
<name>IN_B_0</name></connection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66,-1.5,70.5,-1.5</points>
<intersection>66 2</intersection>
<intersection>70 0</intersection>
<intersection>70.5 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>66,-1.5,66,0.5</points>
<connection>
<GID>245</GID>
<name>OUT_0</name></connection>
<intersection>-1.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>70.5,-20.5,70.5,-1.5</points>
<intersection>-20.5 5</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>70.5,-20.5,71.5,-20.5</points>
<connection>
<GID>37</GID>
<name>IN_B_0</name></connection>
<intersection>70.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-6.5,57.5,-1</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-1,60,-1</points>
<intersection>57.5 0</intersection>
<intersection>60 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>60,-1,60,0.5</points>
<connection>
<GID>244</GID>
<name>OUT_0</name></connection>
<intersection>-1 2</intersection>
<intersection>0.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>60,0.5,61,0.5</points>
<intersection>60 6</intersection>
<intersection>61 10</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>60,-20.5,60,-16.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>-16.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>60,-16.5,61,-16.5</points>
<intersection>60 8</intersection>
<intersection>61 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>61,-16.5,61,0.5</points>
<intersection>-16.5 9</intersection>
<intersection>0.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-6.5,55.5,-1</points>
<connection>
<GID>6</GID>
<name>IN_B_0</name></connection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-1,55.5,-1</points>
<intersection>53 2</intersection>
<intersection>55.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-1,53,1</points>
<connection>
<GID>243</GID>
<name>OUT_0</name></connection>
<intersection>-1 1</intersection>
<intersection>-0.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>53,-0.5,58,-0.5</points>
<intersection>53 2</intersection>
<intersection>58 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>58,-20.5,58,-0.5</points>
<connection>
<GID>36</GID>
<name>IN_B_0</name></connection>
<intersection>-0.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-5.5,44.5,-1.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>44.5,-1.5,46.5,-1.5</points>
<intersection>44.5 0</intersection>
<intersection>46.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>46.5,-1.5,46.5,0.5</points>
<connection>
<GID>242</GID>
<name>OUT_0</name></connection>
<intersection>-1.5 2</intersection>
<intersection>0 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>46.5,0,51.5,0</points>
<intersection>46.5 3</intersection>
<intersection>51.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>51.5,-20.5,51.5,0</points>
<intersection>-20.5 8</intersection>
<intersection>0 4</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>48,-20.5,51.5,-20.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>51.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-8.5,67,-8.5</points>
<connection>
<GID>8</GID>
<name>carry_out</name></connection>
<intersection>60.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>60.5,-9.5,60.5,-8.5</points>
<connection>
<GID>6</GID>
<name>carry_in</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,-8.5,52.5,-8.5</points>
<connection>
<GID>4</GID>
<name>carry_in</name></connection>
<intersection>52.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>52.5,-9.5,52.5,-8.5</points>
<connection>
<GID>6</GID>
<name>carry_out</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-8.5,39.5,-8.5</points>
<connection>
<GID>4</GID>
<name>carry_out</name></connection>
<intersection>36 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-9.5,36,-8.5</points>
<connection>
<GID>2</GID>
<name>carry_in</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-9.5,25.5,-8.5</points>
<intersection>-9.5 2</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-8.5,25.5,-8.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-9.5,28,-9.5</points>
<connection>
<GID>2</GID>
<name>carry_out</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-20.5,46,-15</points>
<connection>
<GID>35</GID>
<name>IN_B_0</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-15,46,-15</points>
<intersection>44.5 2</intersection>
<intersection>46 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>44.5,-15,44.5,-1</points>
<intersection>-15 1</intersection>
<intersection>-1 4</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>42.5,-5.5,42.5,-1</points>
<connection>
<GID>4</GID>
<name>IN_B_0</name></connection>
<intersection>-1 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>41,-1,44.5,-1</points>
<intersection>41 5</intersection>
<intersection>42.5 3</intersection>
<intersection>44.5 2</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>41,-1,41,0.5</points>
<intersection>-1 4</intersection>
<intersection>0.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>40.5,0.5,41,0.5</points>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection>
<intersection>41 5</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-20.5,35.5,-15.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-15.5,36.5,-15.5</points>
<intersection>35.5 0</intersection>
<intersection>36.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>36.5,-15.5,36.5,-6.5</points>
<intersection>-15.5 1</intersection>
<intersection>-6.5 10</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>35.5,-6.5,35.5,0.5</points>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection>
<intersection>-6.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>33,-6.5,36.5,-6.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>35.5 3</intersection>
<intersection>36.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-20.5,31,-16.5</points>
<intersection>-20.5 7</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-16.5,32.5,-16.5</points>
<intersection>31 0</intersection>
<intersection>32.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>32.5,-16.5,32.5,-2</points>
<intersection>-16.5 1</intersection>
<intersection>-2 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>31,-6.5,31,-2</points>
<connection>
<GID>2</GID>
<name>IN_B_0</name></connection>
<intersection>-2 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>28,-2,32.5,-2</points>
<intersection>28 6</intersection>
<intersection>31 4</intersection>
<intersection>32.5 2</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>28,-2,28,0.5</points>
<connection>
<GID>239</GID>
<name>OUT_0</name></connection>
<intersection>-2 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>31,-20.5,33.5,-20.5</points>
<connection>
<GID>34</GID>
<name>IN_B_0</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,-23.5,68.5,-23.5</points>
<connection>
<GID>36</GID>
<name>carry_in</name></connection>
<connection>
<GID>37</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51,-23.5,55,-23.5</points>
<connection>
<GID>36</GID>
<name>carry_out</name></connection>
<connection>
<GID>35</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-23.5,43,-23.5</points>
<connection>
<GID>34</GID>
<name>carry_in</name></connection>
<connection>
<GID>35</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-26.5,26,-12.5</points>
<intersection>-26.5 4</intersection>
<intersection>-12.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>26,-12.5,32,-12.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>26,-26.5,33.5,-26.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-26.5,35.5,-26.5</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-27.5,40,-12</points>
<intersection>-27.5 4</intersection>
<intersection>-12 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>40,-12,43.5,-12</points>
<intersection>40 0</intersection>
<intersection>43.5 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>40,-27.5,48,-27.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>43.5,-12,43.5,-11.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-12 3</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-27.5,50,-27</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47,-27,50,-27</points>
<intersection>47 3</intersection>
<intersection>50 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47,-27,47,-26.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>-27 2</intersection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-28,54,-20</points>
<intersection>-28 3</intersection>
<intersection>-20 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>56.5,-20,56.5,-12.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54,-20,56.5,-20</points>
<intersection>54 0</intersection>
<intersection>56.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>54,-28,62,-28</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-28,64,-27</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>-27 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>59,-27,59,-26.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,-27,64,-27</points>
<intersection>59 1</intersection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-27.5,75,-12.5</points>
<intersection>-27.5 3</intersection>
<intersection>-12.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74.5,-27.5,75,-27.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>71,-12.5,75,-12.5</points>
<intersection>71 5</intersection>
<intersection>75 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>71,-12.5,71,-11.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-12.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-27.5,76.5,-27</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>-27 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>72.5,-27,72.5,-26.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>72.5,-27,76.5,-27</points>
<intersection>72.5 1</intersection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-36.5,36,-33.5</points>
<connection>
<GID>59</GID>
<name>N_in3</name></connection>
<intersection>-33.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>34.5,-33.5,34.5,-30.5</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>-33.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-33.5,36,-33.5</points>
<intersection>34.5 1</intersection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-37,50,-34</points>
<connection>
<GID>61</GID>
<name>N_in3</name></connection>
<intersection>-34 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>49,-34,49,-31.5</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>49,-34,50,-34</points>
<intersection>49 1</intersection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-37,64.5,-34.5</points>
<connection>
<GID>63</GID>
<name>N_in3</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>63,-34.5,63,-32</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,-34.5,64.5,-34.5</points>
<intersection>63 1</intersection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-37,76,-34</points>
<connection>
<GID>65</GID>
<name>N_in3</name></connection>
<intersection>-34 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>75.5,-34,75.5,-31.5</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>75.5,-34,76,-34</points>
<intersection>75.5 1</intersection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-10,16.5,-9.5</points>
<intersection>-10 2</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-9.5,19.5,-9.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-10,16.5,-10</points>
<connection>
<GID>67</GID>
<name>N_in1</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-23.5,27,-10.5</points>
<intersection>-23.5 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-10.5,27,-10.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-23.5,30.5,-23.5</points>
<connection>
<GID>34</GID>
<name>carry_out</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-28.5,21.5,-12</points>
<connection>
<GID>28</GID>
<name>SEL_0</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-28.5,51.5,-28.5</points>
<connection>
<GID>50</GID>
<name>SEL_0</name></connection>
<intersection>21.5 0</intersection>
<intersection>51.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>51.5,-30,51.5,-28.5</points>
<connection>
<GID>51</GID>
<name>SEL_0</name></connection>
<intersection>-30 3</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>51.5,-30,78,-30</points>
<connection>
<GID>52</GID>
<name>SEL_0</name></connection>
<intersection>51.5 2</intersection>
<intersection>78 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78,-30,78,-29.5</points>
<connection>
<GID>53</GID>
<name>SEL_0</name></connection>
<intersection>-30 3</intersection>
<intersection>-29.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>78,-29.5,87.5,-29.5</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<intersection>78 4</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-23.5,79.5,-22.5</points>
<connection>
<GID>256</GID>
<name>OUT_0</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-23.5,79.5,-23.5</points>
<connection>
<GID>37</GID>
<name>carry_in</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-24.1344,0.26646,111.334,-67.8</PageViewport>
<gate>
<ID>195</ID>
<type>FF_GND</type>
<position>31.5,-46.5</position>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>197</ID>
<type>GA_LED</type>
<position>79.5,-47</position>
<input>
<ID>N_in0</ID>98 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>198</ID>
<type>AA_LABEL</type>
<position>15,-23</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>199</ID>
<type>AA_LABEL</type>
<position>27.5,-26</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>200</ID>
<type>AA_LABEL</type>
<position>43,-27</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>AA_LABEL</type>
<position>59.5,-25</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>203</ID>
<type>AA_LABEL</type>
<position>78.5,-42.5</position>
<gparam>LABEL_TEXT Cout</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>205</ID>
<type>AA_LABEL</type>
<position>72,-62.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>206</ID>
<type>AA_LABEL</type>
<position>63,-63.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>207</ID>
<type>AA_LABEL</type>
<position>54.5,-64</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>AA_LABEL</type>
<position>46,-64</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AA_LABEL</type>
<position>38,-63.5</position>
<gparam>LABEL_TEXT S4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>AA_LABEL</type>
<position>46.5,-0.5</position>
<gparam>LABEL_TEXT Carry Save Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>212</ID>
<type>AA_LABEL</type>
<position>22.5,-27</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>213</ID>
<type>AA_LABEL</type>
<position>36.5,-28</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>214</ID>
<type>AA_LABEL</type>
<position>52,-27.5</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>AA_LABEL</type>
<position>68.5,-27.5</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>216</ID>
<type>AA_LABEL</type>
<position>63,-14</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>217</ID>
<type>AA_LABEL</type>
<position>50.5,-14</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>AA_LABEL</type>
<position>38,-14</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_LABEL</type>
<position>25.5,-13.5</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>221</ID>
<type>AA_LABEL</type>
<position>54.5,-66</position>
<gparam>LABEL_TEXT Output</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>AA_LABEL</type>
<position>14,-8.5</position>
<gparam>LABEL_TEXT Inputs</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>224</ID>
<type>AA_LABEL</type>
<position>10,-25</position>
<gparam>LABEL_TEXT Inputs</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>226</ID>
<type>AA_TOGGLE</type>
<position>21.5,-8.5</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>227</ID>
<type>AA_TOGGLE</type>
<position>26,-8</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>228</ID>
<type>AA_TOGGLE</type>
<position>30,-8.5</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_TOGGLE</type>
<position>37.5,-8</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>230</ID>
<type>AA_TOGGLE</type>
<position>41,-8</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>231</ID>
<type>AA_TOGGLE</type>
<position>45,-8.5</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>232</ID>
<type>AA_TOGGLE</type>
<position>50,-8.5</position>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_TOGGLE</type>
<position>54.5,-9</position>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>234</ID>
<type>AA_TOGGLE</type>
<position>59.5,-9</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>235</ID>
<type>AA_TOGGLE</type>
<position>63,-9</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_TOGGLE</type>
<position>66.5,-9</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>237</ID>
<type>AA_TOGGLE</type>
<position>70,-9</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_FULLADDER_1BIT</type>
<position>25,-19</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_B_0</ID>47 </input>
<output>
<ID>OUT_0</ID>59 </output>
<input>
<ID>carry_in</ID>49 </input>
<output>
<ID>carry_out</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_FULLADDER_1BIT</type>
<position>38,-19</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_B_0</ID>50 </input>
<output>
<ID>OUT_0</ID>60 </output>
<input>
<ID>carry_in</ID>52 </input>
<output>
<ID>carry_out</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_FULLADDER_1BIT</type>
<position>51.5,-19.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_B_0</ID>53 </input>
<output>
<ID>OUT_0</ID>68 </output>
<input>
<ID>carry_in</ID>55 </input>
<output>
<ID>carry_out</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_FULLADDER_1BIT</type>
<position>64.5,-19</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_B_0</ID>56 </input>
<output>
<ID>OUT_0</ID>69 </output>
<input>
<ID>carry_in</ID>58 </input>
<output>
<ID>carry_out</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_FULLADDER_1BIT</type>
<position>22.5,-31</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_B_0</ID>65 </input>
<output>
<ID>OUT_0</ID>74 </output>
<input>
<ID>carry_in</ID>82 </input>
<output>
<ID>carry_out</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_FULLADDER_1BIT</type>
<position>36.5,-32</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_B_0</ID>66 </input>
<output>
<ID>OUT_0</ID>76 </output>
<input>
<ID>carry_in</ID>83 </input>
<output>
<ID>carry_out</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_FULLADDER_1BIT</type>
<position>52,-32</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_B_0</ID>67 </input>
<output>
<ID>OUT_0</ID>78 </output>
<input>
<ID>carry_in</ID>84 </input>
<output>
<ID>carry_out</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_FULLADDER_1BIT</type>
<position>67,-32</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_B_0</ID>70 </input>
<output>
<ID>OUT_0</ID>80 </output>
<input>
<ID>carry_in</ID>85 </input>
<output>
<ID>carry_out</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_TOGGLE</type>
<position>17,-26</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_TOGGLE</type>
<position>30.5,-26.5</position>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_TOGGLE</type>
<position>46,-27.5</position>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_TOGGLE</type>
<position>61.5,-26.5</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>156</ID>
<type>AA_FULLADDER_1BIT</type>
<position>27,-43.5</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_B_0</ID>75 </input>
<output>
<ID>OUT_0</ID>88 </output>
<input>
<ID>carry_in</ID>94 </input>
<output>
<ID>carry_out</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_FULLADDER_1BIT</type>
<position>39.5,-43.5</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_B_0</ID>77 </input>
<output>
<ID>OUT_0</ID>89 </output>
<input>
<ID>carry_in</ID>95 </input>
<output>
<ID>carry_out</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>158</ID>
<type>AA_FULLADDER_1BIT</type>
<position>51.5,-43.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_B_0</ID>79 </input>
<output>
<ID>OUT_0</ID>90 </output>
<input>
<ID>carry_in</ID>96 </input>
<output>
<ID>carry_out</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_FULLADDER_1BIT</type>
<position>65,-43.5</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_B_0</ID>81 </input>
<output>
<ID>OUT_0</ID>91 </output>
<input>
<ID>carry_in</ID>97 </input>
<output>
<ID>carry_out</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_LABEL</type>
<position>51.5,-39</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>38.5,-39.5</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>AA_LABEL</type>
<position>26.5,-39</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>AA_LABEL</type>
<position>64.5,-38</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>GA_LED</type>
<position>72,-60.5</position>
<input>
<ID>N_in3</ID>74 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>FF_GND</type>
<position>28,-32.5</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>173</ID>
<type>GA_LED</type>
<position>63,-61</position>
<input>
<ID>N_in3</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>GA_LED</type>
<position>54,-61</position>
<input>
<ID>N_in3</ID>89 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>GA_LED</type>
<position>45.5,-61</position>
<input>
<ID>N_in3</ID>90 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>GA_LED</type>
<position>38.5,-61</position>
<input>
<ID>N_in3</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>21.5,-5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>181</ID>
<type>AA_LABEL</type>
<position>37,-5.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>AA_LABEL</type>
<position>50,-6</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_LABEL</type>
<position>63,-5.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>26,-5.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>AA_LABEL</type>
<position>30,-6</position>
<gparam>LABEL_TEXT C0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>40.5,-5.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>AA_LABEL</type>
<position>54.5,-6</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>188</ID>
<type>AA_LABEL</type>
<position>66,-5.5</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>189</ID>
<type>AA_LABEL</type>
<position>45,-5.5</position>
<gparam>LABEL_TEXT C1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>AA_LABEL</type>
<position>59.5,-5.5</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>191</ID>
<type>AA_LABEL</type>
<position>70,-5.5</position>
<gparam>LABEL_TEXT C3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-16,25.5,-11.5</points>
<intersection>-16 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-11.5,26,-11.5</points>
<intersection>25.5 0</intersection>
<intersection>26 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-16,25.5,-16</points>
<connection>
<GID>120</GID>
<name>IN_B_0</name></connection>
<intersection>25.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>26,-11.5,26,-10</points>
<connection>
<GID>227</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-16,29.5,-12</points>
<intersection>-16 2</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-12,30,-12</points>
<intersection>29.5 0</intersection>
<intersection>30 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-16,29.5,-16</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30,-12,30,-10.5</points>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-14,21,-12</points>
<intersection>-14 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-14,29,-14</points>
<intersection>21 0</intersection>
<intersection>29 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-12,21.5,-12</points>
<intersection>21 0</intersection>
<intersection>21.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>29,-19,29,-14</points>
<connection>
<GID>120</GID>
<name>carry_in</name></connection>
<intersection>-14 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>21.5,-12,21.5,-10.5</points>
<connection>
<GID>226</GID>
<name>OUT_0</name></connection>
<intersection>-12 2</intersection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-16,40.5,-13.5</points>
<intersection>-16 2</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-13.5,41,-13.5</points>
<intersection>40.5 0</intersection>
<intersection>41 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-16,40.5,-16</points>
<connection>
<GID>122</GID>
<name>IN_B_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>41,-13.5,41,-10</points>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection>
<intersection>-13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-16,39,-9.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-9.5,45,-9.5</points>
<intersection>39 0</intersection>
<intersection>45 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>45,-10.5,45,-9.5</points>
<connection>
<GID>231</GID>
<name>OUT_0</name></connection>
<intersection>-9.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-19,43,-10</points>
<intersection>-19 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-19,43,-19</points>
<connection>
<GID>122</GID>
<name>carry_in</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-10,43,-10</points>
<connection>
<GID>229</GID>
<name>OUT_0</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-16.5,54,-11</points>
<intersection>-16.5 2</intersection>
<intersection>-11 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-16.5,54,-16.5</points>
<connection>
<GID>124</GID>
<name>IN_B_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>54,-11,54.5,-11</points>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-16.5,52.5,-11.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-11.5,58,-11.5</points>
<intersection>52.5 0</intersection>
<intersection>58 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>58,-13.5,58,-11.5</points>
<intersection>-13.5 6</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>58,-13.5,59.5,-13.5</points>
<intersection>58 2</intersection>
<intersection>59.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>59.5,-13.5,59.5,-11</points>
<connection>
<GID>234</GID>
<name>OUT_0</name></connection>
<intersection>-13.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-19.5,50,-10.5</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-19.5,55.5,-19.5</points>
<connection>
<GID>124</GID>
<name>carry_in</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-16,66,-11</points>
<intersection>-16 2</intersection>
<intersection>-11 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-16,66,-16</points>
<connection>
<GID>126</GID>
<name>IN_B_0</name></connection>
<intersection>66 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>66,-11,66.5,-11</points>
<connection>
<GID>236</GID>
<name>OUT_0</name></connection>
<intersection>66 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-16,65.5,-12</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-12,70,-12</points>
<intersection>65.5 0</intersection>
<intersection>70 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>70,-12,70,-11</points>
<connection>
<GID>237</GID>
<name>OUT_0</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-19,69,-11.5</points>
<intersection>-19 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-19,69,-19</points>
<connection>
<GID>126</GID>
<name>carry_in</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-11.5,69,-11.5</points>
<intersection>62.5 3</intersection>
<intersection>69 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>62.5,-11.5,62.5,-11</points>
<intersection>-11.5 2</intersection>
<intersection>-11 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>62.5,-11,63,-11</points>
<connection>
<GID>235</GID>
<name>OUT_0</name></connection>
<intersection>62.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-28,23.5,-25</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-25 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>25,-25,25,-22</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-25,25,-25</points>
<intersection>23.5 0</intersection>
<intersection>25 1</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-29,37.5,-25.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>38,-25.5,38,-22</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-25.5,38,-25.5</points>
<intersection>37.5 0</intersection>
<intersection>38 1</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-28,21.5,-26</points>
<connection>
<GID>128</GID>
<name>IN_B_0</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-26,21.5,-26</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-29,35.5,-26.5</points>
<connection>
<GID>130</GID>
<name>IN_B_0</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-26.5,35.5,-26.5</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-29,51,-27.5</points>
<connection>
<GID>132</GID>
<name>IN_B_0</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-27.5,51,-27.5</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-29,53,-25.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>51.5,-25.5,51.5,-22.5</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-25.5,53,-25.5</points>
<intersection>51.5 1</intersection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-29,68,-25.5</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>64.5,-25.5,64.5,-22</points>
<connection>
<GID>126</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-25.5,68,-25.5</points>
<intersection>64.5 1</intersection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-29,66,-26.5</points>
<connection>
<GID>134</GID>
<name>IN_B_0</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-26.5,66,-26.5</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<intersection>66 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-59.5,72,-42</points>
<connection>
<GID>165</GID>
<name>N_in3</name></connection>
<intersection>-42 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>22.5,-42,22.5,-34</points>
<connection>
<GID>128</GID>
<name>OUT_0</name></connection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-42,72,-42</points>
<intersection>22.5 1</intersection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-40.5,26,-36.5</points>
<connection>
<GID>156</GID>
<name>IN_B_0</name></connection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-36.5,26,-36.5</points>
<intersection>18.5 2</intersection>
<intersection>26 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>18.5,-36.5,18.5,-31</points>
<connection>
<GID>128</GID>
<name>carry_out</name></connection>
<intersection>-36.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-40.5,28,-37.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>-37.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>36.5,-37.5,36.5,-35</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28,-37.5,36.5,-37.5</points>
<intersection>28 0</intersection>
<intersection>36.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-40.5,38.5,-36.5</points>
<connection>
<GID>157</GID>
<name>IN_B_0</name></connection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-36.5,38.5,-36.5</points>
<intersection>32.5 2</intersection>
<intersection>38.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>32.5,-36.5,32.5,-32</points>
<connection>
<GID>130</GID>
<name>carry_out</name></connection>
<intersection>-36.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-40.5,40.5,-37.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>-37.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>52,-37.5,52,-35</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-37.5,52,-37.5</points>
<intersection>40.5 0</intersection>
<intersection>52 1</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-40.5,50.5,-32</points>
<connection>
<GID>158</GID>
<name>IN_B_0</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-32,50.5,-32</points>
<connection>
<GID>132</GID>
<name>carry_out</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-40.5,52.5,-37.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>-37.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>67,-37.5,67,-35</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>52.5,-37.5,67,-37.5</points>
<intersection>52.5 0</intersection>
<intersection>67 1</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-40.5,62.5,-32</points>
<intersection>-40.5 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-32,63,-32</points>
<connection>
<GID>134</GID>
<name>carry_out</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-40.5,64,-40.5</points>
<connection>
<GID>159</GID>
<name>IN_B_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-31.5,28,-31</points>
<connection>
<GID>169</GID>
<name>OUT_0</name></connection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-31,28,-31</points>
<connection>
<GID>128</GID>
<name>carry_in</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-24.5,25.5,-23</points>
<intersection>-24.5 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-24.5,40.5,-24.5</points>
<intersection>25.5 0</intersection>
<intersection>40.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-23,25.5,-23</points>
<intersection>21 4</intersection>
<intersection>25.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>40.5,-32,40.5,-24.5</points>
<connection>
<GID>130</GID>
<name>carry_in</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>21,-23,21,-19</points>
<connection>
<GID>120</GID>
<name>carry_out</name></connection>
<intersection>-23 2</intersection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-25.5,41.5,-23</points>
<intersection>-25.5 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-25.5,56,-25.5</points>
<intersection>41.5 0</intersection>
<intersection>56 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-23,41.5,-23</points>
<intersection>34 4</intersection>
<intersection>41.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>56,-32,56,-25.5</points>
<connection>
<GID>132</GID>
<name>carry_in</name></connection>
<intersection>-25.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>34,-23,34,-19</points>
<connection>
<GID>122</GID>
<name>carry_out</name></connection>
<intersection>-23 2</intersection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,-24,71,-24</points>
<intersection>47.5 4</intersection>
<intersection>71 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71,-32,71,-24</points>
<connection>
<GID>134</GID>
<name>carry_in</name></connection>
<intersection>-24 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>47.5,-24,47.5,-19.5</points>
<connection>
<GID>124</GID>
<name>carry_out</name></connection>
<intersection>-24 1</intersection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-40.5,57.5,-19</points>
<intersection>-40.5 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-19,60.5,-19</points>
<connection>
<GID>126</GID>
<name>carry_out</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-40.5,66,-40.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-60,63,-52</points>
<connection>
<GID>173</GID>
<name>N_in3</name></connection>
<intersection>-52 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>27,-52,27,-46.5</points>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27,-52,63,-52</points>
<intersection>27 1</intersection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-60,54,-53.5</points>
<connection>
<GID>176</GID>
<name>N_in3</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>39.5,-53.5,39.5,-46.5</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>39.5,-53.5,54,-53.5</points>
<intersection>39.5 1</intersection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-60,45.5,-48.5</points>
<connection>
<GID>177</GID>
<name>N_in3</name></connection>
<intersection>-48.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>51.5,-48.5,51.5,-46.5</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<intersection>-48.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-48.5,51.5,-48.5</points>
<intersection>45.5 0</intersection>
<intersection>51.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-60,38.5,-51</points>
<connection>
<GID>178</GID>
<name>N_in3</name></connection>
<intersection>-51 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>65,-51,65,-46.5</points>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-51,65,-51</points>
<intersection>38.5 0</intersection>
<intersection>65 1</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-45.5,31.5,-43.5</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-43.5,31.5,-43.5</points>
<connection>
<GID>156</GID>
<name>carry_in</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-41.5,43.5,-41.5</points>
<intersection>23 4</intersection>
<intersection>43.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43.5,-43.5,43.5,-41.5</points>
<connection>
<GID>157</GID>
<name>carry_in</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>23,-43.5,23,-41.5</points>
<connection>
<GID>156</GID>
<name>carry_out</name></connection>
<intersection>-41.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-48,55.5,-48</points>
<intersection>35.5 4</intersection>
<intersection>55.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>55.5,-48,55.5,-43.5</points>
<connection>
<GID>158</GID>
<name>carry_in</name></connection>
<intersection>-48 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>35.5,-48,35.5,-43.5</points>
<connection>
<GID>157</GID>
<name>carry_out</name></connection>
<intersection>-48 1</intersection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,-41.5,69,-41.5</points>
<intersection>47.5 4</intersection>
<intersection>69 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>69,-43.5,69,-41.5</points>
<connection>
<GID>159</GID>
<name>carry_in</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>47.5,-43.5,47.5,-41.5</points>
<connection>
<GID>158</GID>
<name>carry_out</name></connection>
<intersection>-41.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-46,75,-46</points>
<intersection>61 4</intersection>
<intersection>75 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75,-47,75,-46</points>
<intersection>-47 5</intersection>
<intersection>-46 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>61,-46,61,-43.5</points>
<connection>
<GID>159</GID>
<name>carry_out</name></connection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>75,-47,78.5,-47</points>
<connection>
<GID>197</GID>
<name>N_in0</name></connection>
<intersection>75 3</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,33.0808,338.954,-137.227</PageViewport></page 2>
<page 3>
<PageViewport>0,33.0808,338.954,-137.227</PageViewport></page 3>
<page 4>
<PageViewport>0,33.0808,338.954,-137.227</PageViewport></page 4>
<page 5>
<PageViewport>0,33.0808,338.954,-137.227</PageViewport></page 5>
<page 6>
<PageViewport>0,33.0808,338.954,-137.227</PageViewport></page 6>
<page 7>
<PageViewport>0,33.0808,338.954,-137.227</PageViewport></page 7>
<page 8>
<PageViewport>0,33.0808,338.954,-137.227</PageViewport></page 8>
<page 9>
<PageViewport>0,33.0808,338.954,-137.227</PageViewport></page 9></circuit>